//--------------------------------------------------------------------------------------------
// class: Parameterized class
// Description of the class
// class with one parameterized task and one calling task 
//--------------------------------------------------------------------------------------------

class tb#(parameter rx);

//--------------------------------------------------------------------------------------------
// parameterized task 
//--------------------------------------------------------------------------------------------

 task mytask(input bit [rx-1:0]a, input bit [rx-1:0]b);
   bit[rx-1:0] x;
   bit[rx-1:0] y;
   x=a;
   y=b;
   $display("x=%0d,y=%0d,a=%0d,b=%0d",x,y,a,b);
 endtask

//--------------------------------------------------------------------------------------------
// Calling task 
//--------------------------------------------------------------------------------------------
  
 task mytask2;
   bit [rx-1:0]a;
   bit [rx-1:0]b;
   a=8;
   b=11;
   mytask(a,b);
 endtask
  
endclass

//--------------------------------------------------------------------------------------------
// Top module
//--------------------------------------------------------------------------------------------

 module ptask();
  
  tb#(4) p;
  
  initial begin
    p = new();
    p.mytask2;
  end

endmodule
