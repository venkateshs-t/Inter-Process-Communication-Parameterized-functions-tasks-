//--------------------------------------------------------------------------------------------
// wait order in events
//--------------------------------------------------------------------------------------------
module tb;
  event a,b,c;
//--------------------------------------------------------------------------------------------
// process to trigger the events
//--------------------------------------------------------------------------------------------
  initial 
    begin
      #10 -> a;
      #10 -> b;
      #10 -> c;
    end
//--------------------------------------------------------------------------------------------
// wait_order process
//--------------------------------------------------------------------------------------------
  initial 
    begin
      $display("-----------------------------------------------");
      wait_order(a,b,c)
      $display("Events were executed in the correct order");
      else
      $display("Events were not executed in the correct order"); 
      $display("-----------------------------------------------");
    end
  
endmodule
  
      
