//--------------------------------------------------------------------------------------------
//  Merging events
//--------------------------------------------------------------------------------------------
  
module tb;
  event a,b;

  initial 
    begin
      fork
//--------------------------------------------------------------------------------------------
//waiting for event a to trigger 
//--------------------------------------------------------------------------------------------
      begin
        wait(a.triggered);
        $display("@%0d:T1:Wait for event1 is over",$time);
      end
//--------------------------------------------------------------------------------------------
// waiting for event b to trigger
//--------------------------------------------------------------------------------------------
      begin
        wait(b.triggered);
        $display("@%0d:T2:Wait for event2 is over",$time);
      end
//--------------------------------------------------------------------------------------------
// triggering event b
//--------------------------------------------------------------------------------------------
   #30 -> b;
//--------------------------------------------------------------------------------------------
//mergging event b with a 
//--------------------------------------------------------------------------------------------
      begin
        #10 b = a;
      end
    join
  end
  
endmodule
  

